`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2019/02/11 14:41:22
// Design Name: 
// Module Name: InstrDef
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//opcode type
`define U_TYPE  4'b1000
`define J_TYPE  4'b0001
`define B_TYPE  4'b0010
`define L_TYPE  4'b1011
`define S_TYPE  4'b0100
`define I_TYPE  4'b1101
`define R_TYPE  4'b1110

//alu calculate type
`define ALU_ADD 



